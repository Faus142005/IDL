library verilog;
use verilog.vl_types.all;
entity PruebaPrincipal2_vlg_vec_tst is
end PruebaPrincipal2_vlg_vec_tst;
