library verilog;
use verilog.vl_types.all;
entity Registro12_vlg_vec_tst is
end Registro12_vlg_vec_tst;
