library verilog;
use verilog.vl_types.all;
entity PruebaPrincipal_vlg_vec_tst is
end PruebaPrincipal_vlg_vec_tst;
