library verilog;
use verilog.vl_types.all;
entity Registros_vlg_vec_tst is
end Registros_vlg_vec_tst;
