library verilog;
use verilog.vl_types.all;
entity AnalizadorCorte_vlg_vec_tst is
end AnalizadorCorte_vlg_vec_tst;
