library verilog;
use verilog.vl_types.all;
entity Registros_vlg_check_tst is
    port(
        Output          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Registros_vlg_check_tst;
